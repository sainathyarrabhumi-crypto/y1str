package count_package;
int no_of_transactions= 300;
`include "count_trans.sv"
`include "count_gen.sv"
`include "count_wr.sv"
`include "count_wr_mon.sv"
`include "count_ref_model.sv"
`include "count_rd_mon.sv"
`include "count_sb.sv"
`include "count_env.sv"
`include "test.sv"
endpackage
